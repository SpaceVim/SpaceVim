module test1;

reg test;

    test.
test.

mod #(
    .TEST  (1)
) test(
    .port1 (test),
    .
);

mod test(
    .port1 (test),
    .
);

mod
test(
    .port1 (test),
    .
);

 mod #(
    .TEST  (1)
) test(
    .port1 (test),
    .
);

 mod test(
    .port1 (test),
    .port2 (bus[(3-1):0]),
    .port3 (test),
    .in1   (in1),
    .
);

 mod
 test(
    .port1 (test),
    .
);

ola = test.

mod u_mod1 (
    .
);
endmodule

class test2 #(type T=base);

myclass #(type BASE=base) object;
myclass object_with_long_name;
myclass obj;
T typeclass;

object.method(
    .
);

object.atask(.);

object.

object_with_long_name.

obj.

typeclass.

endclass

// vi: set expandtab softtabstop=4 shiftwidth=4:
